// TODO add header

module rr_x_in_tb;

// TODO fill

endmodule;
