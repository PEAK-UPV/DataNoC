// TODO add header

module network_injector_tb;

// TODO fill

endmodule;
