// TODO add header

module switch_2dmesh_vc_tb;

// TODO fill

endmodule;
